module rom0 (
	input  [7:0]  dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [7:0]  dout
);

	RAMB4_S8    RAMA_EXAMPLE (
	    .DO(dout),
	    .ADDR(address),
	    .DI(dinp),
	    .EN(enable),
	    .CLK(clk),
	    .WE(wren),
	    .RST(1'b0)
);

//synthesis attribute INIT_00 of RAMA_EXAMPLE is "BA050E4D494541000000008052004F412020672067206D4D6E704D6F4F6143EB"
//synthesis attribute INIT_01 of RAMA_EXAMPLE is "B304E28817BE0765A20710038804C0E17702E9C1B9902CCD0F4A90CD75E4A835"
//synthesis attribute INIT_02 of RAMA_EXAMPLE is "C613EB74905090FC00C6C7E80B5527E80B03B3E890132CB37490B202E81894BE"
//synthesis attribute INIT_03 of RAMA_EXAMPLE is "9CBE07E814B3902EFF1C90FC2C550BBEFFBE0736BA8B06F613E9137D0480FE03"
//synthesis attribute INIT_04 of RAMA_EXAMPLE is "00843D0F001CCEFC841610FF02569FFFEB468A0710A30014CD10E99059FE01CD"
//synthesis attribute INIT_05 of RAMA_EXAMPLE is "3BFF90F1E48A7300905806C08286DF903E149A90903E20843D00843D0F004BB2"
//synthesis attribute INIT_06 of RAMA_EXAMPLE is "1CCAF64604E53B5E8401FE0001FE0F0DFE0FC3C2E82404468A0F8CE9E95AE888"
//synthesis attribute INIT_07 of RAMA_EXAMPLE is "C3070430C1C60005E80015C3300704810790068904C311EBFE00B9D0C6E92DB9"
//synthesis attribute INIT_08 of RAMA_EXAMPLE is "1E50B404F8050017FD10C7105F478A07C3890A2004070C301B463374C3000607"
//synthesis attribute INIT_09 of RAMA_EXAMPLE is "B458CD8BCD32C358FF530F045A10FF50508E5059FEE8748AB9581F00060404D8"
//synthesis attribute INIT_0A of RAMA_EXAMPLE is "204C0D657420797973500D6464636E632C3267700D306956494F7270202D5820"
//synthesis attribute INIT_0B of RAMA_EXAMPLE is "652020452928726D506165656865206574651869557420754342007520207473"
//synthesis attribute INIT_0C of RAMA_EXAMPLE is "5D6C65395B2020202020206F0404040404030303006E63206E20632020457361"
//synthesis attribute INIT_0D of RAMA_EXAMPLE is "4B47433A61207461366127202020200069003374662046683020202020207364"
//synthesis attribute INIT_0E of RAMA_EXAMPLE is "000000000000000000000000000000000000000000000000000000000074004F"
//synthesis attribute INIT_0F of RAMA_EXAMPLE is "0100000000000000000000000000000000000000000000000000000000000000"

endmodule

module rom1 (
	input  [7:0]  dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [7:0]  dout
);

	RAMB4_S8    RAMB_EXAMPLE (
	    .DO(dout),
	    .ADDR(address),
	    .DI(dinp),
	    .EN(enable),
	    .CLK(clk),
	    .WE(wren),
	    .RST(1'b0)
);

//synthesis attribute INIT_00 of RAMB_EXAMPLE is "0409504C48441200000000004929522F7228616D6F65614F6F4F4F69206F5004"
//synthesis attribute INIT_01 of RAMB_EXAMPLE is "03014704BF0015A1000ECDB4FB2A32C1060EC18100900000EBEA0A0110FA61B9"
//synthesis attribute INIT_02 of RAMB_EXAMPLE is "930E901C90FC1280B4FE8307B2FFBECAB96146700406C690F63506B60500E8D2"
//synthesis attribute INIT_03 of RAMB_EXAMPLE is "E818B30505FF060732FC1480E8FFB2902E02B302902E3008A090068207078B07"
//synthesis attribute INIT_04 of RAMB_EXAMPLE is "3D0F0050C7FC84800FCDCD324DFEE8F0F8050017B90764A000CD75903CEDFC00"
//synthesis attribute INIT_05 of RAMB_EXAMPLE is "4E64903B8490F1C13780F633777224028076729000803C0FB33D0F004DB90084"
//synthesis attribute INIT_06 of RAMB_EXAMPLE is "E8FE75FF8A8490F64644FA3CE9FFF7E9FF00FFFE00887504FFF1E85EC25E56F6"
//synthesis attribute INIT_07 of RAMB_EXAMPLE is "46047204048A04E8000E16072C748AE81102C6E407CF0E46B23CE92A8B5EE820"
//synthesis attribute INIT_08 of RAMB_EXAMPLE is "52C3C3C6E28810BFE6079006F804001707DE042C722C722C74049000FE04C710"
//synthesis attribute INIT_09 of RAMB_EXAMPLE is "515B07010251EA5B3250748A58CD325816C052EF4690C02E515B10B900844A8E"
//synthesis attribute INIT_0A of RAMB_EXAMPLE is "5A410A756E6F656E730A7061696661613120696F302073204252656D73505900"
//synthesis attribute INIT_0B of RAMB_EXAMPLE is "7664743A4E3F656120537467437420746353006C20657270202D0A6E65707220"
//synthesis attribute INIT_0C of RAMB_EXAMPLE is "3175442E202020202020004D7A72614010D4C6AC6C61737361647364743A6568"
//synthesis attribute INIT_0D of RAMB_EXAMPLE is "4A46427466736368314D202020202773725D326C656846305B20202020207364"
//synthesis attribute INIT_0E of RAMB_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000695D4E"
//synthesis attribute INIT_0F of RAMB_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"

endmodule

module rom2 (
	input  [7:0]  dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [7:0]  dout
);

	RAMB4_S8    RAMC_EXAMPLE (
	    .DO(dout),
	    .ADDR(address),
	    .DI(dinp),
	    .EN(enable),
	    .CLK(clk),
	    .WE(wren),
	    .RST(1'b0)
);

//synthesis attribute INIT_00 of RAMC_EXAMPLE is "52BE4F4B4743340000050037432020436F206D61726C535269005274644290AA"
//synthesis attribute INIT_01 of RAMC_EXAMPLE is "7CE8468A0010A307640EFFCBE2F649CBC688010023053DB4E4E275B4A874E400"
//synthesis attribute INIT_02 of RAMC_EXAMPLE is "79FE90FC19807416B9900327902E032A20E803B375388A90858B3003B7BA0533"
//synthesis attribute INIT_03 of RAMC_EXAMPLE is "050002DABA2755278580745F902E070207E2070290F8BFB4FF00C60F1313EB13"
//synthesis attribute INIT_04 of RAMC_EXAMPLE is "0147C00084800F010800025EE88BF0EAE28867BE0015A2C37F0F4E10DF8480B4"
//synthesis attribute INIT_05 of RAMC_EXAMPLE is "248A1CF346903BE87404D85046418C079039301E07A8005374004FA500843D0F"
//synthesis attribute INIT_06 of RAMC_EXAMPLE is "524EC044560F1675048A84804E073B46133C1B010190E488333BFFFFFE015277"
//synthesis attribute INIT_07 of RAMC_EXAMPLE is "04903A04E8C3C6000BE88B1490C0C3000607C33214038BC28480F7C7FE5A00B0"
//synthesis attribute INIT_08 of RAMC_EXAMPLE is "51C346C34604B957E81100C6E28810BF15EBE29010900A90C08A903C37079006"
//synthesis attribute INIT_09 of RAMC_EXAMPLE is "50590EB4B453EB100E90C02E5B09511F8933C3EB009084005059CD07B83616C0"
//synthesis attribute INIT_0A of RAMC_EXAMPLE is "2D280D6E6F746B61650D6A2E7773686D31747243306E72532020746F754910B9"
//synthesis attribute INIT_0B of RAMC_EXAMPLE is "616E69592F2074726500496E3A6E7349653A79697053656D73500D6568756173"
//synthesis attribute INIT_0C of RAMC_EXAMPLE is "3A61202E20202020202065000407040604060306654345656872696E694E6763"
//synthesis attribute INIT_0D of RAMC_EXAMPLE is "4945416C65726143205B2020202020677468317544462E302020202020206541"
//synthesis attribute INIT_0E of RAMC_EXAMPLE is "000000000000000000000000000000000000000000000000000000000078274D"
//synthesis attribute INIT_0F of RAMC_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"

endmodule

module rom3 (
	input  [7:0]  dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [7:0]  dout
);

	RAMB4_S8    RAMD_EXAMPLE (
	    .DO(dout),
	    .ADDR(address),
	    .DI(dinp),
	    .EN(enable),
	    .CLK(clk),
	    .WE(wren),
	    .RST(1'b0)
);

//synthesis attribute INIT_00 of RAMD_EXAMPLE is "E81F4E4A4642010004000076504D54506665497250702020744C6E7072497255"
//synthesis attribute INIT_01 of RAMD_EXAMPLE is "E8F8050767B90014A0893204463309000009FF78E8751690759016FA6110820A"
//synthesis attribute INIT_02 of RAMD_EXAMPLE is "07E52980749048CDEB0847BE02077000B00767900702073D9001BF8BBE039807"
//synthesis attribute INIT_03 of RAMD_EXAMPLE is "F1BAA7BE70E9FFBE0F90FF030457275527E813013503E4077407FF903E069006"
//synthesis attribute INIT_04 of RAMD_EXAMPLE is "1000843D0F0001053CB4B45A520200D74704BF0065A1071025B43C74240F1602"
//synthesis attribute INIT_05 of RAMD_EXAMPLE is "88597375242956901F178E1E3C3C7410903C3C741072AB0052FF00843D0F0048"
//synthesis attribute INIT_06 of RAMD_EXAMPLE is "565E8488FEF7EBC088560FFFCA84FFC28480E984B990842483003C40469304F1"
//synthesis attribute INIT_07 of RAMD_EXAMPLE is "88903CE2C05A0008E80752A29084FE01C7100430A007F4FE0FFE8B2BC4010101"
//synthesis attribute INIT_08 of RAMD_EXAMPLE is "53FF005F478A07C3000607C34605B95716D0C1903C903C9084D22A80E81101C6"
//synthesis attribute INIT_09 of RAMD_EXAMPLE is "C3100E10FF5046CDB49084C359B45304D81E58C2080A0401C35A00B74A8A8A33"
//synthesis attribute INIT_0A of RAMD_EXAMPLE is "540A2E6963202020720A2E652E4063203068790A2E6F654F4D20754342C3CD01"
//synthesis attribute INIT_0B of RAMD_EXAMPLE is "7361780059736561766D206172456D206C1974747520746F7549296D74207469"
//synthesis attribute INIT_0C of RAMD_EXAMPLE is "746620302020202020206400770851BC0081B652633A20676361646178206E20"
//synthesis attribute INIT_0D of RAMD_EXAMPLE is "4844277544657220782020202020206E53343A6120462E302020206820007200"
//synthesis attribute INIT_0E of RAMD_EXAMPLE is "000000000000000000000000000000000000000000000000000000000045504C"
//synthesis attribute INIT_0F of RAMD_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"

endmodule

