module rom(
	input  [31:0] dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [31:0] dout
);

rom3 rom3_inst (
	.dinp(dinp[7:0]),
	.wren(wren),
	.address(address),
	.clk(clk),
	.enable(enable),
	.dout(dout[7:0])
);

rom2 rom2_inst (
	.dinp(dinp[15:8]),
	.wren(wren),
	.address(address),
	.clk(clk),
	.enable(enable),
	.dout(dout[15:8])
);
rom1 rom1_inst (
	.dinp(dinp[23:16]),
	.wren(wren),
	.address(address),
	.clk(clk),
	.enable(enable),
	.dout(dout[23:16])
);
rom0 rom0_inst (
	.dinp(dinp[31:24]),
	.wren(wren),
	.address(address),
	.clk(clk),
	.enable(enable),
	.dout(dout[31:24])
);
endmodule

//-----------------------------------
// これ以降は rom2verilog.c を使って自動生成したものをコピーする
//-----------------------------------

module rom0 (
	input  [7:0]  dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [7:0]  dout
);

	RAMB4_S8    RAMA_EXAMPLE (
	    .DO(dout),
	    .ADDR(address),
	    .DI(dinp),
	    .EN(enable),
	    .CLK(clk),
	    .WE(wren),
	    .RST(1'b0)
);

//synthesis attribute INIT_00 of RAMA_EXAMPLE is "BA050E4D494541000000008052004F412020672067206D4D6E704D6F4F6143EB"
//synthesis attribute INIT_01 of RAMA_EXAMPLE is "B304E288E9BE0665A20610038804C0E17702E9C1B9002CCD0F4A08CD75E4A835"
//synthesis attribute INIT_02 of RAMA_EXAMPLE is "C6E5EB0F005010FC00C6C7E80B95F9E80B03B3E802E52CB30F00B202E81896BE"
//synthesis attribute INIT_03 of RAMA_EXAMPLE is "050002ACBA2595F985800F5F002E060206E2060200F8BF90E5E9E57D0480FE03"
//synthesis attribute INIT_04 of RAMA_EXAMPLE is "0147C00084800F010800025EE88BF0EAE28867BE00E7A2C37F0F4E84DF8480B4"
//synthesis attribute INIT_05 of RAMA_EXAMPLE is "248A83F346273BE80F04D85046418C060039308406A8005374004FA500843D0F"
//synthesis attribute INIT_06 of RAMA_EXAMPLE is "524EC044560F1675048A84804E073B46133C1B010100E488333BFFFFFE015277"
//synthesis attribute INIT_07 of RAMA_EXAMPLE is "04003A04E8C3C6000BE88BE600C0C3000606C332E6038BC28480F7C7FE5A00B0"
//synthesis attribute INIT_08 of RAMA_EXAMPLE is "51C346C34604B957E8E300C6E28810BFE7EBE20010000A00C08A283C37069006"
//synthesis attribute INIT_09 of RAMA_EXAMPLE is "5059E0B4B453EB100E00C02E5B09511F8933C3EB000884005059CD07B83616C0"
//synthesis attribute INIT_0A of RAMA_EXAMPLE is "65616E4D532074490A6E657072205A412E6963202020726D6F65614F6F4F10B9"
//synthesis attribute INIT_0B of RAMA_EXAMPLE is "654345656872696E694E6763616E69592F2074726500496E3A6E7349653A6D6F"
//synthesis attribute INIT_0C of RAMA_EXAMPLE is "44462E3020202020202065413A61202E20202020202065000406040604060306"
//synthesis attribute INIT_0D of RAMA_EXAMPLE is "00000000000000000078274D4945416C65726143205B20202020206774683175"
//synthesis attribute INIT_0E of RAMA_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"
//synthesis attribute INIT_0F of RAMA_EXAMPLE is "5D00000000000000000000000000000000000000000000000000000000000000"

endmodule

module rom1 (
	input  [7:0]  dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [7:0]  dout
);

	RAMB4_S8    RAMB_EXAMPLE (
	    .DO(dout),
	    .ADDR(address),
	    .DI(dinp),
	    .EN(enable),
	    .CLK(clk),
	    .WE(wren),
	    .RST(1'b0)
);

//synthesis attribute INIT_00 of RAMB_EXAMPLE is "040B504C48441200000018004929522F7228616D6F65614F6F4F4F69206F5004"
//synthesis attribute INIT_01 of RAMB_EXAMPLE is "03034704BF00E7A100E0CDB4FB2A32C1060EC18100030000EBEA850110FA61B9"
//synthesis attribute INIT_02 of RAMB_EXAMPLE is "930E001C17FC8480B4FE8106B2FFBECAB96346708506C600F6B506B60500E8D2"
//synthesis attribute INIT_03 of RAMB_EXAMPLE is "C3BAA7BE70E9FFBE0F00FF030457F995F9E8E501B503E408A090068206068B06"
//synthesis attribute INIT_04 of RAMB_EXAMPLE is "1000843D0F0001053CB4B45A520200D74704BF0065A1061025B43C0F240F1602"
//synthesis attribute INIT_05 of RAMB_EXAMPLE is "88590F75248356001F178E1E3C3C74E2123C3C0FE272AB0052FF00843D0F0048"
//synthesis attribute INIT_06 of RAMB_EXAMPLE is "565E8488FEF7EBC088560FFFCA84FFC28480E984B902842483003C40469304F1"
//synthesis attribute INIT_07 of RAMB_EXAMPLE is "88023CE2C05A0008E80652A20584FE01C7E20430A006F4FE0FFE8B2BC4010101"
//synthesis attribute INIT_08 of RAMB_EXAMPLE is "53FF005F478A06C3000606C34605B95716D0C1023C0A3C1984D28480E8E301C6"
//synthesis attribute INIT_09 of RAMB_EXAMPLE is "C3100E10FF5046CDB40D84C359B45304D81E58C208840401C35A00B74A8A8A33"
//synthesis attribute INIT_0A of RAMB_EXAMPLE is "6C53654F4F6E70430D65687561732D286574207979735061726C535269C3CD01"
//synthesis attribute INIT_0B of RAMB_EXAMPLE is "633A20676361646178206E207361780059736561766D206172456D206C196172"
//synthesis attribute INIT_0C of RAMB_EXAMPLE is "20462E30202020682000720074662030202020202020640079DA538E0253B824"
//synthesis attribute INIT_0D of RAMB_EXAMPLE is "00000000000000000045504C4844277544657220782020202020206E53343A61"
//synthesis attribute INIT_0E of RAMB_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"
//synthesis attribute INIT_0F of RAMB_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"

endmodule

module rom2 (
	input  [7:0]  dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [7:0]  dout
);

	RAMB4_S8    RAMC_EXAMPLE (
	    .DO(dout),
	    .ADDR(address),
	    .DI(dinp),
	    .EN(enable),
	    .CLK(clk),
	    .WE(wren),
	    .RST(1'b0)
);

//synthesis attribute INIT_00 of RAMC_EXAMPLE is "54BE4F4B4743340000050068432020436F206D61726C535269005274644290AA"
//synthesis attribute INIT_01 of RAMC_EXAMPLE is "7EE8468A0010A306640EFFCBE2F649CBC688010023853DB4E4E20FB4A874E400"
//synthesis attribute INIT_02 of RAMC_EXAMPLE is "79FE27FC84800F16B90003F9002E032A20E803B30F388A3B858B020389BA0533"
//synthesis attribute INIT_03 of RAMC_EXAMPLE is "BE07E814B3002EFF1C12FC2C950BBEFFBE0736BA8B06F6B4FF00C60FE5E5EBE5"
//synthesis attribute INIT_04 of RAMC_EXAMPLE is "843D0F001CCEFC841610FF02569FFFEB468A0610A300E6CD10E90059FE01CD9C"
//synthesis attribute INIT_05 of RAMC_EXAMPLE is "FF00F1E48A0F00355806C08286DF903E869A00903E20843D00843D0F004BB200"
//synthesis attribute INIT_06 of RAMC_EXAMPLE is "CAF64604E53B5E8401FE0001FE0F0DFE0FC3C2E82485468A0F8CE9E95AE8883B"
//synthesis attribute INIT_07 of RAMC_EXAMPLE is "078230C1C60005E800E7C3308404810690068904C3E3EBFE00B9D0C6E92DB91C"
//synthesis attribute INIT_08 of RAMC_EXAMPLE is "50B404F80500E9FD10C7E25F478A06C3890A20820782308446330FC3000606C3"
//synthesis attribute INIT_09 of RAMC_EXAMPLE is "58CD8BCD32C358FF5384045A10FF50508E5059FEE80F8AB9581F00060404D81E"
//synthesis attribute INIT_0A of RAMC_EXAMPLE is "70204D52496F4F50296D74207469540A756E6F656E730A7250702020745820B4"
//synthesis attribute INIT_0B of RAMC_EXAMPLE is "6E63206E20632020457361652020452928726D50616565686520657465187250"
//synthesis attribute INIT_0C of RAMC_EXAMPLE is "20466830202020202073645D6C65395B2020202020206F040404040403030300"
//synthesis attribute INIT_0D of RAMC_EXAMPLE is "000000000000000074004F4B47433A6120746136612720202020006900337466"
//synthesis attribute INIT_0E of RAMC_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"
//synthesis attribute INIT_0F of RAMC_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"

endmodule

module rom3 (
	input  [7:0]  dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [7:0]  dout
);

	RAMB4_S8    RAMD_EXAMPLE (
	    .DO(dout),
	    .ADDR(address),
	    .DI(dinp),
	    .EN(enable),
	    .CLK(clk),
	    .WE(wren),
	    .RST(1'b0)
);

//synthesis attribute INIT_00 of RAMD_EXAMPLE is "E81F4E4A4642010004000009504D54506665497250702020744C6E7072497255"
//synthesis attribute INIT_01 of RAMD_EXAMPLE is "E8F8050667B900E6A0893204463309000009FF78E80F1690750016FA6110821E"
//synthesis attribute INIT_02 of RAMD_EXAMPLE is "06E584800F0048CDEB0849BE02067200B0076900060207840001BF8DBE036107"
//synthesis attribute INIT_03 of RAMD_EXAMPLE is "18B30505FF060630FC8480E8FFB2002E02B302002E0290067406FF903E069006"
//synthesis attribute INIT_04 of RAMD_EXAMPLE is "0F0050C7FC84800FCDCD324DFEE8F0F80500E9B90664A000CD750E3CEBFC00E8"
//synthesis attribute INIT_05 of RAMD_EXAMPLE is "641A3B8400F1C18480F63377722402800F721C00803C0FB33D0F004DB900843D"
//synthesis attribute INIT_06 of RAMD_EXAMPLE is "FE75FF8A8490F64644FA3CE9FFF7E9FF00FFFE00880F04FFF1E85EC25E56F64E"
//synthesis attribute INIT_07 of RAMD_EXAMPLE is "040F04048A04E8000E16062C0F8AE8E302C6E406CF0E46B23CE92A8B5EE820E8"
//synthesis attribute INIT_08 of RAMD_EXAMPLE is "C3C3C6E28810BFE6069006F80400E906DE042C0F2C0F2C0F040000FE04C7E246"
//synthesis attribute INIT_09 of RAMD_EXAMPLE is "5B06010251EA5B32500F8A58CD325816C052EF4600C02E515B10B900844A8E52"
//synthesis attribute INIT_0A of RAMD_EXAMPLE is "6D752020426920007520207473204C0D6E6F746B61650D67206D4D6E70590051"
//synthesis attribute INIT_0B of RAMD_EXAMPLE is "61737361647364743A65687664743A4E3F656120537467437420746353006720"
//synthesis attribute INIT_0C of RAMD_EXAMPLE is "6846305B202020202073643175442E202020202020004D7C74634212D6C8AE6C"
//synthesis attribute INIT_0D of RAMD_EXAMPLE is "0000000000000000695D4E4A46427466736368314D202020202773725D326C65"
//synthesis attribute INIT_0E of RAMD_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"
//synthesis attribute INIT_0F of RAMD_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"

endmodule

