module rom0 (
	input  [7:0]  dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [7:0]  dout
);

	RAMB4_S8    RAMA_EXAMPLE (
	    .DO(dout),
	    .ADDR(address),
	    .DI(dinp),
	    .EN(enable),
	    .CLK(clk),
	    .WE(wren),
	    .RST(1'b0)
);

//synthesis attribute INIT_00 of RAMA_EXAMPLE is "BA050E20202F49000000008052004F412020672067206D4D6E704D6F4F6143EB"
//synthesis attribute INIT_01 of RAMA_EXAMPLE is "03014704BF002FA10028CDB4FB2A32C1060EC181CB902CCD0F4A90CD75E4A835"
//synthesis attribute INIT_02 of RAMA_EXAMPLE is "930E901C90FC1280B4FE8307B2FFBECAB96146700406C690F63506B60500E8D2"
//synthesis attribute INIT_03 of RAMA_EXAMPLE is "E818B30505FF060732FC1480E8FFB2902E02B302902E3608A090068207078B07"
//synthesis attribute INIT_04 of RAMA_EXAMPLE is "3D0F0050C7FC84800FCDCD324DFEE8F0F8050031B90764A000CD75903CEDFC00"
//synthesis attribute INIT_05 of RAMA_EXAMPLE is "4E64903B8490F1C13780F633777224028076729000803C0FB33D0F004DB90084"
//synthesis attribute INIT_06 of RAMA_EXAMPLE is "E8FE75FF8A8490F64644FA3CE9FFF7E9FF00FFFE00887504FFF1E85EC25E56F6"
//synthesis attribute INIT_07 of RAMA_EXAMPLE is "46047204048A04E8000E16072C748AE82B02C6E407CF0E46B23CE92A8B5EE820"
//synthesis attribute INIT_08 of RAMA_EXAMPLE is "52C3C3C6E28810BFE6079006F804003107DE042C722C722C74049000FE04C72A"
//synthesis attribute INIT_09 of RAMA_EXAMPLE is "515B07010251EA5B3250748A58CD325816C052EF4690C02E515B10B900844A8E"
//synthesis attribute INIT_0A of RAMA_EXAMPLE is "280D6E6F746B61650D6A2E7773686D313820696F302073204252656D73505900"
//synthesis attribute INIT_0B of RAMA_EXAMPLE is "6E69592F2074726500496E3A6E7349653A79697053656D73500D65687561732D"
//synthesis attribute INIT_0C of RAMA_EXAMPLE is "31202020202020207063000407040604060306654345656872696E694E676361"
//synthesis attribute INIT_0D of RAMA_EXAMPLE is "202020206C74003174662030305B20202020006E6169535D54202B3A53207253"
//synthesis attribute INIT_0E of RAMA_EXAMPLE is "000000000000000000000000000000000000000000000078736368314D202020"
//synthesis attribute INIT_0F of RAMA_EXAMPLE is "5A00000000000000000000000000000000000000000000000000000000000000"

endmodule

module rom1 (
	input  [7:0]  dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [7:0]  dout
);

	RAMB4_S8    RAMB_EXAMPLE (
	    .DO(dout),
	    .ADDR(address),
	    .DI(dinp),
	    .EN(enable),
	    .CLK(clk),
	    .WE(wren),
	    .RST(1'b0)
);

//synthesis attribute INIT_00 of RAMB_EXAMPLE is "040A202050340000000000004929522F7228616D6F65614F6F4F4F69206F5004"
//synthesis attribute INIT_01 of RAMB_EXAMPLE is "7CE8468A0010A307640EFFCBE2F649CBC688010000900000EBEA0A0110FA61B9"
//synthesis attribute INIT_02 of RAMB_EXAMPLE is "79FE90FC19807416B9900341902E032A20E803B375388A90858B3603BDBA0533"
//synthesis attribute INIT_03 of RAMB_EXAMPLE is "050002E0BA2755418580745F902E070207E2070290F8BFB4FF00C60F2D2DEB2D"
//synthesis attribute INIT_04 of RAMB_EXAMPLE is "0147C00084800F010800025EE88BF0EAE28867BE002FA2C37F0F4E10DF8480B4"
//synthesis attribute INIT_05 of RAMB_EXAMPLE is "248A1CF346903BE87404D85046418C079039301E07A8005374004FA500843D0F"
//synthesis attribute INIT_06 of RAMB_EXAMPLE is "524EC044560F1675048A84804E073B46133C1B010190E488333BFFFFFE015277"
//synthesis attribute INIT_07 of RAMB_EXAMPLE is "04903A04E8C3C6000BE88B2E90C0C3000607C3322E038BC28480F7C7FE5A00B0"
//synthesis attribute INIT_08 of RAMB_EXAMPLE is "51C346C34604B957E82B00C6E28810BF2FEBE29010900A90C08A903C37079006"
//synthesis attribute INIT_09 of RAMB_EXAMPLE is "505928B4B453EB100E90C02E5B09511F8933C3EB009084005059CD07B83616C0"
//synthesis attribute INIT_0A of RAMB_EXAMPLE is "0A2E6963202020720A2E652E4063203030747243306E72532020746F754910B9"
//synthesis attribute INIT_0B of RAMB_EXAMPLE is "61780059736561766D206172456D206C1974747520746F7549296D7420746954"
//synthesis attribute INIT_0C of RAMB_EXAMPLE is "5B20202020202020796E00782252E801A5B758633A20676361646178206E2073"
//synthesis attribute INIT_0D of RAMB_EXAMPLE is "202020206F6F5D306C653030302020202020296F7A7455524F4D533344726955"
//synthesis attribute INIT_0E of RAMB_EXAMPLE is "000000000000000000000000000000000000000000000045726143205B202020"
//synthesis attribute INIT_0F of RAMB_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"

endmodule

module rom2 (
	input  [7:0]  dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [7:0]  dout
);

	RAMB4_S8    RAMC_EXAMPLE (
	    .DO(dout),
	    .ADDR(address),
	    .DI(dinp),
	    .EN(enable),
	    .CLK(clk),
	    .WE(wren),
	    .RST(1'b0)
);

//synthesis attribute INIT_00 of RAMC_EXAMPLE is "53BE20204456100000050037432020436F206D61726C535269005274644290AA"
//synthesis attribute INIT_01 of RAMC_EXAMPLE is "E8F8050767B9002EA0893204463309000009FF7824053DB4E4E275B4A874E400"
//synthesis attribute INIT_02 of RAMC_EXAMPLE is "07E52980749048CDEB0847BE02077000B00767900702073D9001BF8BBE039E07"
//synthesis attribute INIT_03 of RAMC_EXAMPLE is "F7BAA7BE70E9FFBE0F90FF030457415541E82D013503E4077407FF903E069006"
//synthesis attribute INIT_04 of RAMC_EXAMPLE is "1000843D0F0001053CB4B45A520200D74704BF0065A1071025B43C74240F1602"
//synthesis attribute INIT_05 of RAMC_EXAMPLE is "88597375242956901F178E1E3C3C742A903C3C742A72AB0052FF00843D0F0048"
//synthesis attribute INIT_06 of RAMC_EXAMPLE is "565E8488FEF7EBC088560FFFCA84FFC28480E984B990842483003C40469304F1"
//synthesis attribute INIT_07 of RAMC_EXAMPLE is "88903CE2C05A0008E80752A29084FE01C72A0430A007F4FE0FFE8B2BC4010101"
//synthesis attribute INIT_08 of RAMC_EXAMPLE is "53FF005F478A07C3000607C34605B95716D0C1903C903C9084D22A80E82B01C6"
//synthesis attribute INIT_09 of RAMC_EXAMPLE is "C3100E10FF5046CDB49084C359B45304D81E58C2080A0401C35A00B74A8A8A33"
//synthesis attribute INIT_0A of RAMC_EXAMPLE is "0D657420797973500D6464636E632C323068790A2E6F654F4D20754342C3CD01"
//synthesis attribute INIT_0B of RAMC_EXAMPLE is "20452928726D506165656865206574651869557420754342007520207473204C"
//synthesis attribute INIT_0C of RAMC_EXAMPLE is "202020202020200054790404040404030303006E63206E206320204573616520"
//synthesis attribute INIT_0D of RAMC_EXAMPLE is "20202020637220307544302E3020202020202569695542453A5355203A6F4D42"
//synthesis attribute INIT_0E of RAMC_EXAMPLE is "0000000000000000000000000000000000000000000074006572207820202020"
//synthesis attribute INIT_0F of RAMC_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"

endmodule

module rom3 (
	input  [7:0]  dinp,
	input         wren,
	input  [8:0]  address,
	input         clk,
	input         enable,
	output [7:0]  dout
);

	RAMB4_S8    RAMD_EXAMPLE (
	    .DO(dout),
	    .ADDR(address),
	    .DI(dinp),
	    .EN(enable),
	    .CLK(clk),
	    .WE(wren),
	    .RST(1'b0)
);

//synthesis attribute INIT_00 of RAMD_EXAMPLE is "E81F20205550010004000076504D54506665497250702020744C6E7072497255"
//synthesis attribute INIT_01 of RAMD_EXAMPLE is "04E28831BE0765A20710038804C0E17702E9C1B9E8751690759016FA61108203"
//synthesis attribute INIT_02 of RAMD_EXAMPLE is "2DEB74905090FC00C6C7E8155541E81503B3E8902D2CB37490B202E81894BEB3"
//synthesis attribute INIT_03 of RAMD_EXAMPLE is "BE07E814B3902EFF1C90FC2C5515BEFFBE0736BA8B06F62DE92D7D0480FE03C6"
//synthesis attribute INIT_04 of RAMD_EXAMPLE is "843D0F001CCEFC841610FF02569FFFEB468A0710A3002ECD10E99059FE01CD9C"
//synthesis attribute INIT_05 of RAMD_EXAMPLE is "FF90F1E48A7300905806C08286DF903E149A90903E20843D00843D0F004BB200"
//synthesis attribute INIT_06 of RAMD_EXAMPLE is "CAF64604E53B5E8401FE0001FE0F0DFE0FC3C2E82404468A0F8CE9E95AE8883B"
//synthesis attribute INIT_07 of RAMD_EXAMPLE is "070430C1C60005E8002FC3300704810790068904C32BEBFE00B9D0C6E92DB91C"
//synthesis attribute INIT_08 of RAMD_EXAMPLE is "50B404F8050031FD10C72A5F478A07C3890A2004070C301B463374C3000607C3"
//synthesis attribute INIT_09 of RAMD_EXAMPLE is "58CD8BCD32C358FF530F045A10FF50508E5059FEE8748AB9581F00060404D81E"
//synthesis attribute INIT_0A of RAMD_EXAMPLE is "0A756E6F656E730A706169666161312D3267700D306956494F7270202D5820B4"
//synthesis attribute INIT_0B of RAMD_EXAMPLE is "743A4E3F656120537467437420746353006C20657270202D0A6E657072205A41"
//synthesis attribute INIT_0C of RAMD_EXAMPLE is "202020202020206520537B73624111D5C7AD6C61737361647364743A65687664"
//synthesis attribute INIT_0D of RAMD_EXAMPLE is "202020006F50303A6120312E30202020202028746C2000483444424D3272203A"
//synthesis attribute INIT_0E of RAMD_EXAMPLE is "00000000000000000000000000000000000000000000695D7461366120202020"
//synthesis attribute INIT_0F of RAMD_EXAMPLE is "0000000000000000000000000000000000000000000000000000000000000000"

endmodule

